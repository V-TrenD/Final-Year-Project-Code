--
entity KeypadEncoderl is
	port(
		
	);
end KeypadEncoderl;